-------------------------------
-- Gera um pulso se o botÃ£o estiver apertado. SÃ³ comparar
-- se b_out vale '1' num IF para utilizar.
----------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.all;
----------------------------------
ENTITY roleta IS
	PORT (b_in: IN STD_LOGIC;
		  clk: IN STD_LOGIC;
		  r_num: OUT INTEGER);
END ENTITY;
----------------------------------
ARCHITECTURE roleta OF roleta IS
	SIGNAL s_b_in: STD_LOGIC;
	
BEGIN
	PROCESS(clk)
		VARIABLE temp: INTEGER RANGE 1 TO 9;
	BEGIN
		IF (rising_edge(clk)) THEN
			IF(temp >= 9) THEN
				temp := 1;
			ELSE
				temp := temp + 1;
			END IF;
		END IF;

		IF(b_in = '1') THEN
			r_num <= temp;
		END IF;
	END PROCESS;
END ARCHITECTURE;